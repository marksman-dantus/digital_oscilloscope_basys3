library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity char_rom_minimal is
    Port (
        clk         : in  STD_LOGIC;
        char_addr   : in  STD_LOGIC_VECTOR(4 downto 0); -- 32 characters
        row         : in  STD_LOGIC_VECTOR(3 downto 0); -- 16 rows
        col         : in  STD_LOGIC_VECTOR(2 downto 0); -- 8 columns
        char_pixel  : out STD_LOGIC
    );
end char_rom_minimal;

architecture Behavioral of char_rom_minimal is
    -- Define font as a 3D array of std_logic for direct bit access
    type font_array is array (0 to 31, 0 to 15, 0 to 7) of STD_LOGIC;
    constant font : font_array := (
        -- T
        ( ("1","1","1","1","1","1","1","1"), ("1","1","1","1","1","1","1","1"), ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"),
          ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"),
          ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"),
          ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0") ),
        -- r
        ( ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0"),
          ("0","0","0","0","0","0","0","0"), ("0","1","1","1","1","1","0","0"), ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","0","0","0"),
          ("0","1","1","0","0","0","0","0"), ("0","1","1","0","0","0","0","0"), ("0","1","1","0","0","0","0","0"), ("0","1","1","0","0","0","0","0"),
          ("0","1","1","0","0","0","0","0"), ("0","1","1","0","0","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0") ),
        -- i
        ( ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"),
          ("0","0","0","0","0","0","0","0"), ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"),
          ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"),
          ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0") ),
        -- g
        ( ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0"),
          ("0","0","0","0","0","0","0","0"), ("0","0","1","1","1","1","1","0"), ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"),
          ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"),
          ("0","1","1","0","0","1","1","0"), ("0","0","1","1","1","1","1","0"), ("0","0","0","0","0","1","1","0"), ("0","0","1","1","1","1","0","0") ),
        -- :
        ( ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0"),
          ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0"),
          ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","1","1","0","0","0"),
          ("0","0","0","1","1","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0") ),
        -- Space
        ( others => ("0","0","0","0","0","0","0","0") ),
        -- 0
        ( ("0","0","1","1","1","1","0","0"), ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"),
          ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"),
          ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"),
          ("0","1","1","0","0","1","1","0"), ("0","0","1","1","1","1","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0") ),
        -- 1
        ( ("0","0","0","1","1","0","0","0"), ("0","0","1","1","1","0","0","0"), ("0","1","1","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"),
          ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"),
          ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"),
          ("0","0","0","1","1","0","0","0"), ("0","0","1","1","1","1","1","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0") ),
        -- 2
        ( ("0","0","1","1","1","1","0","0"), ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"),
          ("0","0","0","0","0","1","1","0"), ("0","0","0","0","0","1","1","0"), ("0","0","0","0","1","1","0","0"), ("0","0","0","1","1","0","0","0"),
          ("0","0","1","1","0","0","0","0"), ("0","1","1","0","0","0","0","0"), ("0","1","1","0","0","0","0","0"), ("0","1","1","0","0","0","0","0"),
          ("0","1","1","0","0","0","0","0"), ("0","1","1","1","1","1","1","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0") ),
        -- 5
        ( ("0","1","1","1","1","1","1","0"), ("0","1","1","0","0","0","0","0"), ("0","1","1","0","0","0","0","0"), ("0","1","1","0","0","0","0","0"),
          ("0","1","1","0","0","0","0","0"), ("0","1","1","1","1","1","0","0"), ("0","1","1","0","0","1","1","0"), ("0","0","0","0","0","1","1","0"),
          ("0","0","0","0","0","1","1","0"), ("0","0","0","0","0","1","1","0"), ("0","0","0","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"),
          ("0","1","1","0","0","1","1","0"), ("0","0","1","1","1","1","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0") ),
        -- V
        ( ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"),
          ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"),
          ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"), ("0","0","1","1","1","1","0","0"),
          ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0") ),
        -- /
        ( ("0","0","0","0","0","1","1","0"), ("0","0","0","0","0","1","1","0"), ("0","0","0","0","1","1","0","0"), ("0","0","0","0","1","1","0","0"),
          ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"), ("0","0","1","1","0","0","0","0"),
          ("0","0","1","1","0","0","0","0"), ("0","1","1","0","0","0","0","0"), ("0","1","1","0","0","0","0","0"), ("0","1","1","0","0","0","0","0"),
          ("0","1","1","0","0","0","0","0"), ("0","1","1","0","0","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0") ),
        -- d
        ( ("0","0","0","0","0","1","1","0"), ("0","0","0","0","0","1","1","0"), ("0","0","0","0","0","1","1","0"), ("0","0","0","0","0","1","1","0"),
          ("0","0","0","0","0","1","1","0"), ("0","0","1","1","1","1","1","0"), ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"),
          ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"),
          ("0","1","1","0","0","1","1","0"), ("0","0","1","1","1","1","1","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0") ),
        -- ?
        ( ("0","0","1","1","1","1","0","0"), ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"), ("0","0","0","0","0","1","1","0"),
          ("0","0","0","0","0","1","1","0"), ("0","0","0","0","1","1","0","0"), ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"),
          ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0"),
          ("0","0","0","1","1","0","0","0"), ("0","0","0","1","1","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0") ),
        -- P
        ( ("0","1","1","1","1","1","0","0"), ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"),
          ("0","1","1","0","0","1","1","0"), ("0","1","1","0","0","1","1","0"), ("0","1","1","1","1","1","0","0"), ("0","1","1","0","0","0","0","0"),
          ("0","1","1","0","0","0","0","0"), ("0","1","1","0","0","0","0","0"), ("0","1","1","0","0","0","0","0"), ("0","1","1","0","0","0","0","0"),
          ("0","1","1","0","0","0","0","0"), ("0","1","1","0","0","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0") ),
        -- .
        ( ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0"),
          ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0"),
          ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","1","1","0","0","0"),
          ("0","0","0","1","1","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0"), ("0","0","0","0","0","0","0","0") ),
        others => (others => ("0","0","0","0","0","0","0","0"))
    );
begin
    process(clk)
        variable row_idx : integer range 0 to 15;
        variable char_idx : integer range 0 to 31;
        variable col_idx : integer range 0 to 7;
    begin
        if rising_edge(clk) then
            row_idx := to_integer(unsigned(row));
            char_idx := to_integer(unsigned(char_addr));
            col_idx := 7 - to_integer(unsigned(col)); -- Flip column for correct display
            if row_idx < 16 and char_idx < 32 and col_idx < 8 then
                char_pixel <= font(char_idx, row_idx, col_idx);
            else
                char_pixel <= '0';
            end if;
        end if;
    end process;
end Behavioral;