library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity character_rom is
    Port ( 
        clk         : in  STD_LOGIC;
        char_code   : in  STD_LOGIC_VECTOR(7 downto 0);   -- ASCII kodu
        char_x      : in  STD_LOGIC_VECTOR(2 downto 0);   -- 0-7 karakter içi x pozisyonu
        char_y      : in  STD_LOGIC_VECTOR(3 downto 0);   -- 0-15 karakter içi y pozisyonu
        char_pixel  : out STD_LOGIC                       -- Karakter pikseli (1=açık, 0=kapalı)
    );
end character_rom;

architecture Behavioral of character_rom is
    -- 8x16 karakterler için ROM
    type char_rom_t is array (0 to 127, 0 to 15) of std_logic_vector(7 downto 0);
    
    -- Temel ASCII karakterleri içeren ROM. Sadece belli başlı işaretler ve sayılar
    -- Gerçek uygulamada daha fazla karakter eklenebilir
    constant CHAR_ROM : char_rom_t := (
        -- ASCII 32: SPACE
        32 => (
            "00000000", -- 0
            "00000000", -- 1
            "00000000", -- 2
            "00000000", -- 3
            "00000000", -- 4
            "00000000", -- 5
            "00000000", -- 6
            "00000000", -- 7
            "00000000", -- 8
            "00000000", -- 9
            "00000000", -- 10
            "00000000", -- 11
            "00000000", -- 12
            "00000000", -- 13
            "00000000", -- 14
            "00000000"  -- 15
        ),
        -- ASCII 48-57: 0-9
        -- 0
        48 => (
            "00000000", -- 0
            "00111100", -- 1
            "01100110", -- 2
            "01100110", -- 3
            "01100110", -- 4
            "01100110", -- 5
            "01100110", -- 6
            "01100110", -- 7
            "01100110", -- 8
            "01100110", -- 9
            "01100110", -- 10
            "01100110", -- 11
            "00111100", -- 12
            "00000000", -- 13
            "00000000", -- 14
            "00000000"  -- 15
        ),
        -- 1
        49 => (
            "00000000", -- 0
            "00011000", -- 1
            "00111000", -- 2
            "01111000", -- 3
            "00011000", -- 4
            "00011000", -- 5
            "00011000", -- 6
            "00011000", -- 7
            "00011000", -- 8
            "00011000", -- 9
            "00011000", -- 10
            "00011000", -- 11
            "01111110", -- 12
            "00000000", -- 13
            "00000000", -- 14
            "00000000"  -- 15
        ),
        -- 2
        50 => (
            "00000000", -- 0
            "00111100", -- 1
            "01100110", -- 2
            "00000110", -- 3
            "00000110", -- 4
            "00001100", -- 5
            "00011000", -- 6
            "00110000", -- 7
            "01100000", -- 8
            "01100000", -- 9
            "01100000", -- 10
            "01100000", -- 11
            "01111110", -- 12
            "00000000", -- 13
            "00000000", -- 14
            "00000000"  -- 15
        ),
        -- 3
        51 => (
            "00000000", -- 0
            "00111100", -- 1
            "01100110", -- 2
            "00000110", -- 3
            "00000110", -- 4
            "00000110", -- 5
            "00111100", -- 6
            "00000110", -- 7
            "00000110", -- 8
            "00000110", -- 9
            "00000110", -- 10
            "01100110", -- 11
            "00111100", -- 12
            "00000000", -- 13
            "00000000", -- 14
            "00000000"  -- 15
        ),
        -- 4
        52 => (
            "00000000", -- 0
            "00000110", -- 1
            "00001110", -- 2
            "00011110", -- 3
            "00110110", -- 4
            "01100110", -- 5
            "01100110", -- 6
            "01111110", -- 7
            "00000110", -- 8
            "00000110", -- 9
            "00000110", -- 10
            "00000110", -- 11
            "00000110", -- 12
            "00000000", -- 13
            "00000000", -- 14
            "00000000"  -- 15
        ),
        -- 5
        53 => (
            "00000000", -- 0
            "01111110", -- 1
            "01100000", -- 2
            "01100000", -- 3
            "01100000", -- 4
            "01100000", -- 5
            "01111100", -- 6
            "00000110", -- 7
            "00000110", -- 8
            "00000110", -- 9
            "00000110", -- 10
            "01100110", -- 11
            "00111100", -- 12
            "00000000", -- 13
            "00000000", -- 14
            "00000000"  -- 15
        ),
        -- 6
        54 => (
            "00000000", -- 0
            "00111100", -- 1
            "01100110", -- 2
            "01100000", -- 3
            "01100000", -- 4
            "01100000", -- 5
            "01111100", -- 6
            "01100110", -- 7
            "01100110", -- 8
            "01100110", -- 9
            "01100110", -- 10
            "01100110", -- 11
            "00111100", -- 12
            "00000000", -- 13
            "00000000", -- 14
            "00000000"  -- 15
        ),
        -- 7
        55 => (
            "00000000", -- 0
            "01111110", -- 1
            "00000110", -- 2
            "00000110", -- 3
            "00000110", -- 4
            "00001100", -- 5
            "00011000", -- 6
            "00110000", -- 7
            "00110000", -- 8
            "00110000", -- 9
            "00110000", -- 10
            "00110000", -- 11
            "00110000", -- 12
            "00000000", -- 13
            "00000000", -- 14
            "00000000"  -- 15
        ),
        -- 8
        56 => (
            "00000000", -- 0
            "00111100", -- 1
            "01100110", -- 2
            "01100110", -- 3
            "01100110", -- 4
            "01100110", -- 5
            "00111100", -- 6
            "01100110", -- 7
            "01100110", -- 8
            "01100110", -- 9
            "01100110", -- 10
            "01100110", -- 11
            "00111100", -- 12
            "00000000", -- 13
            "00000000", -- 14
            "00000000"  -- 15
        ),
        -- 9
        57 => (
            "00000000", -- 0
            "00111100", -- 1
            "01100110", -- 2
            "01100110", -- 3
            "01100110", -- 4
            "01100110", -- 5
            "00111110", -- 6
            "00000110", -- 7
            "00000110", -- 8
            "00000110", -- 9
            "00000110", -- 10
            "01100110", -- 11
            "00111100", -- 12
            "00000000", -- 13
            "00000000", -- 14
            "00000000"  -- 15
        ),
        -- ASCII 46: dot (.)
        46 => (
            "00000000", -- 0
            "00000000", -- 1
            "00000000", -- 2
            "00000000", -- 3
            "00000000", -- 4
            "00000000", -- 5
            "00000000", -- 6
            "00000000", -- 7
            "00000000", -- 8
            "00000000", -- 9
            "00000000", -- 10
            "00011000", -- 11
            "00011000", -- 12
            "00000000", -- 13
            "00000000", -- 14
            "00000000"  -- 15
        ),
        -- ASCII 86: V
        86 => (
            "00000000", -- 0
            "01100110", -- 1
            "01100110", -- 2
            "01100110", -- 3
            "01100110", -- 4
            "01100110", -- 5
            "01100110", -- 6
            "01100110", -- 7
            "01100110", -- 8
            "01100110", -- 9
            "01100110", -- 10
            "00111100", -- 11
            "00011000", -- 12
            "00000000", -- 13
            "00000000", -- 14
            "00000000"  -- 15
        ),
        -- ASCII 84: T
        84 => (
            "00000000", -- 0
            "01111110", -- 1
            "00011000", -- 2
            "00011000", -- 3
            "00011000", -- 4
            "00011000", -- 5
            "00011000", -- 6
            "00011000", -- 7
            "00011000", -- 8
            "00011000", -- 9
            "00011000", -- 10
            "00011000", -- 11
            "00011000", -- 12
            "00000000", -- 13
            "00000000", -- 14
            "00000000"  -- 15
        ),
        -- ASCII 47: / (slash)
        47 => (
            "00000000", -- 0
            "00000110", -- 1
            "00000110", -- 2
            "00001100", -- 3
            "00001100", -- 4
            "00011000", -- 5
            "00011000", -- 6
            "00110000", -- 7
            "00110000", -- 8
            "01100000", -- 9
            "01100000", -- 10
            "01000000", -- 11
            "01000000", -- 12
            "00000000", -- 13
            "00000000", -- 14
            "00000000"  -- 15
        ),
        -- ASCII 100: d
        100 => (
            "00000000", -- 0
            "00000110", -- 1
            "00000110", -- 2
            "00000110", -- 3
            "00000110", -- 4
            "00111110", -- 5
            "01100110", -- 6
            "01100110", -- 7
            "01100110", -- 8
            "01100110", -- 9
            "01100110", -- 10
            "01100110", -- 11
            "00111110", -- 12
            "00000000", -- 13
            "00000000", -- 14
            "00000000"  -- 15
        ),
        -- ASCII 105: i
        105 => (
            "00000000", -- 0
            "00011000", -- 1
            "00011000", -- 2
            "00000000", -- 3
            "00000000", -- 4
            "00111000", -- 5
            "00011000", -- 6
            "00011000", -- 7
            "00011000", -- 8
            "00011000", -- 9
            "00011000", -- 10
            "00011000", -- 11
            "01111110", -- 12
            "00000000", -- 13
            "00000000", -- 14
            "00000000"  -- 15
        ),
        -- ASCII 118: v
        118 => (
            "00000000", -- 0
            "00000000", -- 1
            "00000000", -- 2
            "00000000", -- 3
            "00000000", -- 4
            "01100110", -- 5
            "01100110", -- 6
            "01100110", -- 7
            "01100110", -- 8
            "01100110", -- 9
            "01100110", -- 10
            "00111100", -- 11
            "00011000", -- 12
            "00000000", -- 13
            "00000000", -- 14
            "00000000"  -- 15
        ),
        -- ASCII 109: m
        109 => (
            "00000000", -- 0
            "00000000", -- 1
            "00000000", -- 2
            "00000000", -- 3
            "00000000", -- 4
            "01100011", -- 5
            "01110111", -- 6
            "01111111", -- 7
            "01101011", -- 8
            "01100011", -- 9
            "01100011", -- 10
            "01100011", -- 11
            "01100011", -- 12
            "00000000", -- 13
            "00000000", -- 14
            "00000000"  -- 15
        ),
        -- ASCII 115: s
        115 => (
            "00000000", -- 0
            "00000000", -- 1
            "00000000", -- 2
            "00000000", -- 3
            "00000000", -- 4
            "00111100", -- 5
            "01100110", -- 6
            "01100000", -- 7
            "00111100", -- 8
            "00000110", -- 9
            "00000110", -- 10
            "01100110", -- 11
            "00111100", -- 12
            "00000000", -- 13
            "00000000", -- 14
            "00000000"  -- 15
        ),
        -- ASCII 83: S
        83 => (
            "00000000", -- 0
            "00111100", -- 1
            "01100110", -- 2
            "01100110", -- 3
            "01100000", -- 4
            "00110000", -- 5
            "00011100", -- 6
            "00000110", -- 7
            "00000110", -- 8
            "00000110", -- 9
            "01100110", -- 10
            "01100110", -- 11
            "00111100", -- 12
            "00000000", -- 13
            "00000000", -- 14
            "00000000"  -- 15
        ),
        -- ASCII 77: M
        77 => (
            "00000000", -- 0
            "01100011", -- 1
            "01110111", -- 2
            "01111111", -- 3
            "01111111", -- 4
            "01101011", -- 5
            "01100011", -- 6
            "01100011", -- 7
            "01100011", -- 8
            "01100011", -- 9
            "01100011", -- 10
            "01100011", -- 11
            "01100011", -- 12
            "00000000", -- 13
            "00000000", -- 14
            "00000000"  -- 15
        ),
        -- ASCII 117: u
        117 => (
            "00000000", -- 0
            "00000000", -- 1
            "00000000", -- 2
            "00000000", -- 3
            "00000000", -- 4
            "01100110", -- 5
            "01100110", -- 6
            "01100110", -- 7
            "01100110", -- 8
            "01100110", -- 9
            "01100110", -- 10
            "01100110", -- 11
            "00111110", -- 12
            "00000000", -- 13
            "00000000", -- 14
            "00000000"  -- 15
        ),
        -- ASCII 58: : (colon)
        58 => (
            "00000000", -- 0
            "00000000", -- 1
            "00000000", -- 2
            "00011000", -- 3
            "00011000", -- 4
            "00000000", -- 5
            "00000000", -- 6
            "00000000", -- 7
            "00000000", -- 8
            "00011000", -- 9
            "00011000", -- 10
            "00000000", -- 11
            "00000000", -- 12
            "00000000", -- 13
            "00000000", -- 14
            "00000000"  -- 15
        ),
        -- ASCII 66: B
        66 => (
            "00000000", -- 0
            "01111100", -- 1
            "01100110", -- 2
            "01100110", -- 3
            "01100110", -- 4
            "01100110", -- 5
            "01111100", -- 6
            "01100110", -- 7
            "01100110", -- 8
            "01100110", -- 9
            "01100110", -- 10
            "01100110", -- 11
            "01111100", -- 12
            "00000000", -- 13
            "00000000", -- 14
            "00000000"  -- 15
        ),
        -- Diğer karakterler için varsayılan (boşluk)
        others => (others => "00000000")
    );
    
    signal rom_addr : integer range 0 to 127;
    signal rom_data : std_logic_vector(7 downto 0);
    signal col_addr : integer range 0 to 7;
    
begin
    -- ASCII kodu 0-127 arasında sınırla
    rom_addr <= to_integer(unsigned(char_code)) when unsigned(char_code) < 128 else 32;
    
    -- Sütun adresi 0-7 arasında
    col_addr <= to_integer(unsigned(char_x));
    
    -- ROM'dan veri alma
    rom_data <= CHAR_ROM(rom_addr, to_integer(unsigned(char_y)));
    
    -- İstenen piksel değerini çıkışa gönder
    char_pixel <= rom_data(7 - col_addr);
    
end Behavioral;